`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    02:03:00 09/16/2014 
// Design Name: 
// Module Name:    segClkDevider 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//��Ƶ����clk_divƵ��ΪԭƵ�ʵ�20000��֮һ���ߵ�ƽ��λ
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module segClkDevider(
input clk,
    input rst,
    output reg clk_div
    );
     
 localparam constantNumber = 10000;
 reg [31:0] count;
 
always @ (posedge(clk), posedge(rst))
begin
    if (rst == 1'b1)
        count <= 32'b0;
    else if (count == constantNumber - 1)
        count <= 32'b0;               
    else
        count <= count + 1;
end

always @ (posedge(clk), posedge(rst))
begin
    if (rst == 1'b1)
        clk_div <= 1'b0;
    else if (count == constantNumber - 1)
        clk_div <= ~clk_div;
    else
        clk_div <= clk_div;
end
endmodule